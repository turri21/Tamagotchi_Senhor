// Build ID Verilog Module
`define BUILD_DATE "20250305"
`define BUILD_HASH "FEEDC0DE"
